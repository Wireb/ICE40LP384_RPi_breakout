-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 1 2022 22:16:29

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "spi_shifter" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of spi_shifter
entity spi_shifter is
port (
    SPI_SS : in std_logic;
    SPI_SDO : out std_logic;
    SPI_SDI : in std_logic;
    LED : out std_logic;
    SPI_SCK : in std_logic);
end spi_shifter;

-- Architecture of spi_shifter
-- View name is \INTERFACE\
architecture \INTERFACE\ of spi_shifter is

signal \N__2548\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2448\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2394\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2367\ : std_logic;
signal \N__2364\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2313\ : std_logic;
signal \N__2310\ : std_logic;
signal \N__2307\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2271\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2256\ : std_logic;
signal \N__2253\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2211\ : std_logic;
signal \N__2208\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2196\ : std_logic;
signal \N__2193\ : std_logic;
signal \N__2190\ : std_logic;
signal \N__2187\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2181\ : std_logic;
signal \N__2178\ : std_logic;
signal \N__2175\ : std_logic;
signal \N__2172\ : std_logic;
signal \N__2169\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2163\ : std_logic;
signal \N__2160\ : std_logic;
signal \N__2157\ : std_logic;
signal \N__2154\ : std_logic;
signal \N__2151\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2145\ : std_logic;
signal \N__2142\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2136\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2127\ : std_logic;
signal \N__2124\ : std_logic;
signal \N__2121\ : std_logic;
signal \N__2118\ : std_logic;
signal \N__2115\ : std_logic;
signal \N__2112\ : std_logic;
signal \N__2109\ : std_logic;
signal \N__2106\ : std_logic;
signal \N__2103\ : std_logic;
signal \N__2100\ : std_logic;
signal \N__2097\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2088\ : std_logic;
signal \N__2085\ : std_logic;
signal \N__2082\ : std_logic;
signal \N__2079\ : std_logic;
signal \N__2076\ : std_logic;
signal \N__2073\ : std_logic;
signal \N__2070\ : std_logic;
signal \N__2067\ : std_logic;
signal \N__2064\ : std_logic;
signal \N__2061\ : std_logic;
signal \N__2058\ : std_logic;
signal \N__2055\ : std_logic;
signal \N__2052\ : std_logic;
signal \N__2049\ : std_logic;
signal \N__2046\ : std_logic;
signal \N__2043\ : std_logic;
signal \N__2040\ : std_logic;
signal \N__2037\ : std_logic;
signal \N__2034\ : std_logic;
signal \N__2031\ : std_logic;
signal \N__2028\ : std_logic;
signal \N__2025\ : std_logic;
signal \N__2022\ : std_logic;
signal \N__2019\ : std_logic;
signal \N__2016\ : std_logic;
signal \N__2013\ : std_logic;
signal \N__2010\ : std_logic;
signal \N__2007\ : std_logic;
signal \N__2004\ : std_logic;
signal \N__2001\ : std_logic;
signal \N__1998\ : std_logic;
signal \N__1995\ : std_logic;
signal \N__1992\ : std_logic;
signal \N__1989\ : std_logic;
signal \N__1986\ : std_logic;
signal \N__1983\ : std_logic;
signal \N__1980\ : std_logic;
signal \N__1977\ : std_logic;
signal \N__1974\ : std_logic;
signal \N__1971\ : std_logic;
signal \N__1968\ : std_logic;
signal \N__1965\ : std_logic;
signal \N__1962\ : std_logic;
signal \N__1959\ : std_logic;
signal \N__1956\ : std_logic;
signal \N__1953\ : std_logic;
signal \N__1950\ : std_logic;
signal \N__1947\ : std_logic;
signal \N__1944\ : std_logic;
signal \N__1941\ : std_logic;
signal \N__1938\ : std_logic;
signal \N__1935\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1929\ : std_logic;
signal \N__1926\ : std_logic;
signal \N__1923\ : std_logic;
signal \N__1920\ : std_logic;
signal \N__1917\ : std_logic;
signal \N__1914\ : std_logic;
signal \N__1911\ : std_logic;
signal \N__1908\ : std_logic;
signal \N__1905\ : std_logic;
signal \N__1902\ : std_logic;
signal \N__1899\ : std_logic;
signal \N__1896\ : std_logic;
signal \N__1893\ : std_logic;
signal \N__1890\ : std_logic;
signal \N__1887\ : std_logic;
signal \N__1884\ : std_logic;
signal \N__1881\ : std_logic;
signal \N__1878\ : std_logic;
signal \N__1875\ : std_logic;
signal \N__1872\ : std_logic;
signal \N__1869\ : std_logic;
signal \N__1866\ : std_logic;
signal \N__1863\ : std_logic;
signal \N__1860\ : std_logic;
signal \N__1857\ : std_logic;
signal \N__1854\ : std_logic;
signal \N__1851\ : std_logic;
signal \N__1848\ : std_logic;
signal \N__1845\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1839\ : std_logic;
signal \N__1836\ : std_logic;
signal \N__1833\ : std_logic;
signal \N__1830\ : std_logic;
signal \N__1827\ : std_logic;
signal \N__1824\ : std_logic;
signal \N__1821\ : std_logic;
signal \N__1818\ : std_logic;
signal \N__1815\ : std_logic;
signal \N__1812\ : std_logic;
signal \N__1809\ : std_logic;
signal \N__1806\ : std_logic;
signal \N__1803\ : std_logic;
signal \N__1800\ : std_logic;
signal \N__1797\ : std_logic;
signal \N__1794\ : std_logic;
signal \N__1791\ : std_logic;
signal \N__1788\ : std_logic;
signal \N__1785\ : std_logic;
signal \N__1782\ : std_logic;
signal \N__1779\ : std_logic;
signal \N__1776\ : std_logic;
signal \N__1773\ : std_logic;
signal \N__1770\ : std_logic;
signal \N__1767\ : std_logic;
signal \N__1764\ : std_logic;
signal \N__1761\ : std_logic;
signal \N__1758\ : std_logic;
signal \N__1755\ : std_logic;
signal \N__1752\ : std_logic;
signal \N__1749\ : std_logic;
signal \N__1746\ : std_logic;
signal \N__1743\ : std_logic;
signal \N__1740\ : std_logic;
signal \N__1737\ : std_logic;
signal \N__1734\ : std_logic;
signal \N__1731\ : std_logic;
signal \N__1728\ : std_logic;
signal \N__1725\ : std_logic;
signal \N__1722\ : std_logic;
signal \N__1719\ : std_logic;
signal \N__1716\ : std_logic;
signal \N__1713\ : std_logic;
signal \N__1710\ : std_logic;
signal \N__1707\ : std_logic;
signal \N__1704\ : std_logic;
signal \N__1701\ : std_logic;
signal \N__1698\ : std_logic;
signal \N__1695\ : std_logic;
signal \N__1692\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1686\ : std_logic;
signal \N__1683\ : std_logic;
signal \N__1680\ : std_logic;
signal \N__1677\ : std_logic;
signal \N__1674\ : std_logic;
signal \N__1671\ : std_logic;
signal \N__1668\ : std_logic;
signal \N__1665\ : std_logic;
signal \N__1662\ : std_logic;
signal \N__1659\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1655\ : std_logic;
signal \N__1654\ : std_logic;
signal \N__1653\ : std_logic;
signal \N__1652\ : std_logic;
signal \N__1651\ : std_logic;
signal \N__1650\ : std_logic;
signal \N__1649\ : std_logic;
signal \N__1648\ : std_logic;
signal \N__1647\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1644\ : std_logic;
signal \N__1643\ : std_logic;
signal \N__1642\ : std_logic;
signal \N__1641\ : std_logic;
signal \N__1640\ : std_logic;
signal \N__1605\ : std_logic;
signal \N__1602\ : std_logic;
signal \N__1599\ : std_logic;
signal \N__1596\ : std_logic;
signal \N__1593\ : std_logic;
signal \N__1590\ : std_logic;
signal \N__1587\ : std_logic;
signal \SPI_SCK_c_g\ : std_logic;
signal \SPI_SCK_ibuf_gb_io_gb_input\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \SPI_SDO_c\ : std_logic;
signal \shift_regZ0Z_119\ : std_logic;
signal \shift_regZ0Z_118\ : std_logic;
signal \shift_regZ0Z_117\ : std_logic;
signal \shift_regZ0Z_116\ : std_logic;
signal \shift_regZ0Z_115\ : std_logic;
signal \INVSPI_SDOZ0C_net\ : std_logic;
signal \shift_regZ0Z_20\ : std_logic;
signal \shift_regZ0Z_21\ : std_logic;
signal \shift_regZ0Z_22\ : std_logic;
signal \shift_regZ0Z_23\ : std_logic;
signal \shift_regZ0Z_24\ : std_logic;
signal \shift_regZ0Z_25\ : std_logic;
signal \shift_regZ0Z_26\ : std_logic;
signal \INVshift_reg_20C_net\ : std_logic;
signal \shift_regZ0Z_27\ : std_logic;
signal \shift_regZ0Z_28\ : std_logic;
signal \shift_regZ0Z_29\ : std_logic;
signal \shift_regZ0Z_30\ : std_logic;
signal \shift_regZ0Z_31\ : std_logic;
signal \shift_regZ0Z_32\ : std_logic;
signal \shift_regZ0Z_33\ : std_logic;
signal \shift_regZ0Z_34\ : std_logic;
signal \INVshift_reg_28C_net\ : std_logic;
signal \shift_regZ0Z_35\ : std_logic;
signal \shift_regZ0Z_36\ : std_logic;
signal \shift_regZ0Z_37\ : std_logic;
signal \shift_regZ0Z_38\ : std_logic;
signal \shift_regZ0Z_39\ : std_logic;
signal \shift_regZ0Z_40\ : std_logic;
signal \shift_regZ0Z_41\ : std_logic;
signal \shift_regZ0Z_42\ : std_logic;
signal \INVshift_reg_36C_net\ : std_logic;
signal \shift_regZ0Z_98\ : std_logic;
signal \shift_regZ0Z_99\ : std_logic;
signal \shift_regZ0Z_100\ : std_logic;
signal \INVshift_reg_98C_net\ : std_logic;
signal \shift_regZ0Z_114\ : std_logic;
signal \shift_regZ0Z_101\ : std_logic;
signal \shift_regZ0Z_102\ : std_logic;
signal \shift_regZ0Z_110\ : std_logic;
signal \shift_regZ0Z_111\ : std_logic;
signal \shift_regZ0Z_112\ : std_logic;
signal \shift_regZ0Z_113\ : std_logic;
signal \INVshift_reg_114C_net\ : std_logic;
signal \shift_regZ0Z_108\ : std_logic;
signal \shift_regZ0Z_109\ : std_logic;
signal \shift_regZ0Z_103\ : std_logic;
signal \shift_regZ0Z_104\ : std_logic;
signal \shift_regZ0Z_105\ : std_logic;
signal \shift_regZ0Z_106\ : std_logic;
signal \shift_regZ0Z_107\ : std_logic;
signal \shift_regZ0Z_18\ : std_logic;
signal \shift_regZ0Z_19\ : std_logic;
signal \INVshift_reg_108C_net\ : std_logic;
signal \shift_regZ0Z_43\ : std_logic;
signal \shift_regZ0Z_44\ : std_logic;
signal \shift_regZ0Z_45\ : std_logic;
signal \shift_regZ0Z_46\ : std_logic;
signal \shift_regZ0Z_47\ : std_logic;
signal \shift_regZ0Z_48\ : std_logic;
signal \shift_regZ0Z_49\ : std_logic;
signal \shift_regZ0Z_50\ : std_logic;
signal \INVshift_reg_44C_net\ : std_logic;
signal \shift_regZ0Z_96\ : std_logic;
signal \shift_regZ0Z_97\ : std_logic;
signal \shift_regZ0Z_6\ : std_logic;
signal \INVshift_reg_96C_net\ : std_logic;
signal \shift_regZ0Z_91\ : std_logic;
signal \shift_regZ0Z_92\ : std_logic;
signal \shift_regZ0Z_93\ : std_logic;
signal \shift_regZ0Z_94\ : std_logic;
signal \shift_regZ0Z_95\ : std_logic;
signal \shift_regZ0Z_7\ : std_logic;
signal \shift_regZ0Z_8\ : std_logic;
signal \INVshift_reg_9C_net\ : std_logic;
signal \shift_regZ0Z_9\ : std_logic;
signal \shift_regZ0Z_10\ : std_logic;
signal \shift_regZ0Z_11\ : std_logic;
signal \shift_regZ0Z_12\ : std_logic;
signal \shift_regZ0Z_13\ : std_logic;
signal \shift_regZ0Z_14\ : std_logic;
signal \shift_regZ0Z_15\ : std_logic;
signal \shift_regZ0Z_16\ : std_logic;
signal \shift_regZ0Z_17\ : std_logic;
signal \INVshift_reg_10C_net\ : std_logic;
signal \shift_regZ0Z_60\ : std_logic;
signal \shift_regZ0Z_61\ : std_logic;
signal \shift_regZ0Z_62\ : std_logic;
signal \shift_regZ0Z_63\ : std_logic;
signal \shift_regZ0Z_64\ : std_logic;
signal \shift_regZ0Z_65\ : std_logic;
signal \shift_regZ0Z_66\ : std_logic;
signal \INVshift_reg_60C_net\ : std_logic;
signal \shift_regZ0Z_51\ : std_logic;
signal \shift_regZ0Z_52\ : std_logic;
signal \shift_regZ0Z_53\ : std_logic;
signal \shift_regZ0Z_54\ : std_logic;
signal \shift_regZ0Z_55\ : std_logic;
signal \shift_regZ0Z_56\ : std_logic;
signal \shift_regZ0Z_57\ : std_logic;
signal \shift_regZ0Z_58\ : std_logic;
signal \shift_regZ0Z_59\ : std_logic;
signal \INVshift_reg_52C_net\ : std_logic;
signal \SPI_SDI_c\ : std_logic;
signal \shift_regZ0Z_0\ : std_logic;
signal \shift_regZ0Z_1\ : std_logic;
signal \shift_regZ0Z_2\ : std_logic;
signal \shift_regZ0Z_3\ : std_logic;
signal \shift_regZ0Z_4\ : std_logic;
signal \shift_regZ0Z_5\ : std_logic;
signal \INVshift_reg_0C_net\ : std_logic;
signal \shift_regZ0Z_90\ : std_logic;
signal \shift_regZ0Z_84\ : std_logic;
signal \shift_regZ0Z_85\ : std_logic;
signal \shift_regZ0Z_86\ : std_logic;
signal \shift_regZ0Z_87\ : std_logic;
signal \shift_regZ0Z_88\ : std_logic;
signal \shift_regZ0Z_89\ : std_logic;
signal \INVshift_reg_90C_net\ : std_logic;
signal \shift_regZ0Z_76\ : std_logic;
signal \shift_regZ0Z_77\ : std_logic;
signal \shift_regZ0Z_78\ : std_logic;
signal \shift_regZ0Z_79\ : std_logic;
signal \shift_regZ0Z_80\ : std_logic;
signal \shift_regZ0Z_81\ : std_logic;
signal \shift_regZ0Z_82\ : std_logic;
signal \shift_regZ0Z_83\ : std_logic;
signal \INVshift_reg_76C_net\ : std_logic;
signal \shift_regZ0Z_67\ : std_logic;
signal \shift_regZ0Z_68\ : std_logic;
signal \shift_regZ0Z_69\ : std_logic;
signal \shift_regZ0Z_70\ : std_logic;
signal \shift_regZ0Z_71\ : std_logic;
signal \shift_regZ0Z_72\ : std_logic;
signal \shift_regZ0Z_73\ : std_logic;
signal \shift_regZ0Z_74\ : std_logic;
signal \shift_regZ0Z_75\ : std_logic;
signal \INVshift_reg_68C_net\ : std_logic;
signal \LED_c_i_g\ : std_logic;
signal \LED_c\ : std_logic;
signal \LED_c_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \SPI_SDO_wire\ : std_logic;
signal \SPI_SDI_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \SPI_SS_wire\ : std_logic;
signal \SPI_SCK_wire\ : std_logic;

begin
    SPI_SDO <= \SPI_SDO_wire\;
    \SPI_SDI_wire\ <= SPI_SDI;
    LED <= \LED_wire\;
    \SPI_SS_wire\ <= SPI_SS;
    \SPI_SCK_wire\ <= SPI_SCK;

    \SPI_SDO_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2548\,
            DIN => \N__2547\,
            DOUT => \N__2546\,
            PACKAGEPIN => \SPI_SDO_wire\
        );

    \SPI_SDO_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2548\,
            PADOUT => \N__2547\,
            PADIN => \N__2546\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1692\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SPI_SDI_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2539\,
            DIN => \N__2538\,
            DOUT => \N__2537\,
            PACKAGEPIN => \SPI_SDI_wire\
        );

    \SPI_SDI_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2539\,
            PADOUT => \N__2538\,
            PADIN => \N__2537\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SPI_SDI_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2530\,
            DIN => \N__2529\,
            DOUT => \N__2528\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2530\,
            PADOUT => \N__2529\,
            PADIN => \N__2528\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2388\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SPI_SS_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2521\,
            DIN => \N__2520\,
            DOUT => \N__2519\,
            PACKAGEPIN => \SPI_SS_wire\
        );

    \SPI_SS_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2521\,
            PADOUT => \N__2520\,
            PADIN => \N__2519\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \LED_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SPI_SCK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2512\,
            DIN => \N__2511\,
            DOUT => \N__2510\,
            PACKAGEPIN => \SPI_SCK_wire\
        );

    \SPI_SCK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2512\,
            PADOUT => \N__2511\,
            PADIN => \N__2510\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SPI_SCK_ibuf_gb_io_gb_input\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__451\ : InMux
    port map (
            O => \N__2493\,
            I => \N__2490\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2490\,
            I => \shift_regZ0Z_68\
        );

    \I__449\ : InMux
    port map (
            O => \N__2487\,
            I => \N__2484\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__2484\,
            I => \shift_regZ0Z_69\
        );

    \I__447\ : InMux
    port map (
            O => \N__2481\,
            I => \N__2478\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__2478\,
            I => \shift_regZ0Z_70\
        );

    \I__445\ : InMux
    port map (
            O => \N__2475\,
            I => \N__2472\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2472\,
            I => \shift_regZ0Z_71\
        );

    \I__443\ : InMux
    port map (
            O => \N__2469\,
            I => \N__2466\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2466\,
            I => \shift_regZ0Z_72\
        );

    \I__441\ : InMux
    port map (
            O => \N__2463\,
            I => \N__2460\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2460\,
            I => \shift_regZ0Z_73\
        );

    \I__439\ : InMux
    port map (
            O => \N__2457\,
            I => \N__2454\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2454\,
            I => \shift_regZ0Z_74\
        );

    \I__437\ : InMux
    port map (
            O => \N__2451\,
            I => \N__2448\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2448\,
            I => \shift_regZ0Z_75\
        );

    \I__435\ : CEMux
    port map (
            O => \N__2445\,
            I => \N__2394\
        );

    \I__434\ : CEMux
    port map (
            O => \N__2444\,
            I => \N__2394\
        );

    \I__433\ : CEMux
    port map (
            O => \N__2443\,
            I => \N__2394\
        );

    \I__432\ : CEMux
    port map (
            O => \N__2442\,
            I => \N__2394\
        );

    \I__431\ : CEMux
    port map (
            O => \N__2441\,
            I => \N__2394\
        );

    \I__430\ : CEMux
    port map (
            O => \N__2440\,
            I => \N__2394\
        );

    \I__429\ : CEMux
    port map (
            O => \N__2439\,
            I => \N__2394\
        );

    \I__428\ : CEMux
    port map (
            O => \N__2438\,
            I => \N__2394\
        );

    \I__427\ : CEMux
    port map (
            O => \N__2437\,
            I => \N__2394\
        );

    \I__426\ : CEMux
    port map (
            O => \N__2436\,
            I => \N__2394\
        );

    \I__425\ : CEMux
    port map (
            O => \N__2435\,
            I => \N__2394\
        );

    \I__424\ : CEMux
    port map (
            O => \N__2434\,
            I => \N__2394\
        );

    \I__423\ : CEMux
    port map (
            O => \N__2433\,
            I => \N__2394\
        );

    \I__422\ : CEMux
    port map (
            O => \N__2432\,
            I => \N__2394\
        );

    \I__421\ : CEMux
    port map (
            O => \N__2431\,
            I => \N__2394\
        );

    \I__420\ : CEMux
    port map (
            O => \N__2430\,
            I => \N__2394\
        );

    \I__419\ : CEMux
    port map (
            O => \N__2429\,
            I => \N__2394\
        );

    \I__418\ : GlobalMux
    port map (
            O => \N__2394\,
            I => \N__2391\
        );

    \I__417\ : gio2CtrlBuf
    port map (
            O => \N__2391\,
            I => \LED_c_i_g\
        );

    \I__416\ : IoInMux
    port map (
            O => \N__2388\,
            I => \N__2384\
        );

    \I__415\ : InMux
    port map (
            O => \N__2387\,
            I => \N__2381\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2384\,
            I => \N__2378\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2381\,
            I => \N__2375\
        );

    \I__412\ : Odrv4
    port map (
            O => \N__2378\,
            I => \LED_c\
        );

    \I__411\ : Odrv4
    port map (
            O => \N__2375\,
            I => \LED_c\
        );

    \I__410\ : IoInMux
    port map (
            O => \N__2370\,
            I => \N__2367\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2367\,
            I => \N__2364\
        );

    \I__408\ : IoSpan4Mux
    port map (
            O => \N__2364\,
            I => \N__2361\
        );

    \I__407\ : Span4Mux_s1_h
    port map (
            O => \N__2361\,
            I => \N__2358\
        );

    \I__406\ : Span4Mux_h
    port map (
            O => \N__2358\,
            I => \N__2355\
        );

    \I__405\ : Odrv4
    port map (
            O => \N__2355\,
            I => \LED_c_i\
        );

    \I__404\ : InMux
    port map (
            O => \N__2352\,
            I => \N__2349\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2349\,
            I => \shift_regZ0Z_76\
        );

    \I__402\ : InMux
    port map (
            O => \N__2346\,
            I => \N__2343\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2343\,
            I => \shift_regZ0Z_77\
        );

    \I__400\ : InMux
    port map (
            O => \N__2340\,
            I => \N__2337\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2337\,
            I => \shift_regZ0Z_78\
        );

    \I__398\ : InMux
    port map (
            O => \N__2334\,
            I => \N__2331\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2331\,
            I => \shift_regZ0Z_79\
        );

    \I__396\ : InMux
    port map (
            O => \N__2328\,
            I => \N__2325\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2325\,
            I => \shift_regZ0Z_80\
        );

    \I__394\ : InMux
    port map (
            O => \N__2322\,
            I => \N__2319\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2319\,
            I => \shift_regZ0Z_81\
        );

    \I__392\ : InMux
    port map (
            O => \N__2316\,
            I => \N__2313\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2313\,
            I => \shift_regZ0Z_82\
        );

    \I__390\ : InMux
    port map (
            O => \N__2310\,
            I => \N__2307\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2307\,
            I => \shift_regZ0Z_83\
        );

    \I__388\ : InMux
    port map (
            O => \N__2304\,
            I => \N__2301\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2301\,
            I => \shift_regZ0Z_67\
        );

    \I__386\ : InMux
    port map (
            O => \N__2298\,
            I => \N__2295\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2295\,
            I => \shift_regZ0Z_3\
        );

    \I__384\ : InMux
    port map (
            O => \N__2292\,
            I => \N__2289\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2289\,
            I => \shift_regZ0Z_4\
        );

    \I__382\ : InMux
    port map (
            O => \N__2286\,
            I => \N__2283\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2283\,
            I => \shift_regZ0Z_5\
        );

    \I__380\ : InMux
    port map (
            O => \N__2280\,
            I => \N__2277\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2277\,
            I => \shift_regZ0Z_90\
        );

    \I__378\ : InMux
    port map (
            O => \N__2274\,
            I => \N__2271\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2271\,
            I => \shift_regZ0Z_84\
        );

    \I__376\ : InMux
    port map (
            O => \N__2268\,
            I => \N__2265\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2265\,
            I => \shift_regZ0Z_85\
        );

    \I__374\ : InMux
    port map (
            O => \N__2262\,
            I => \N__2259\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2259\,
            I => \shift_regZ0Z_86\
        );

    \I__372\ : InMux
    port map (
            O => \N__2256\,
            I => \N__2253\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2253\,
            I => \shift_regZ0Z_87\
        );

    \I__370\ : InMux
    port map (
            O => \N__2250\,
            I => \N__2247\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2247\,
            I => \shift_regZ0Z_88\
        );

    \I__368\ : InMux
    port map (
            O => \N__2244\,
            I => \N__2241\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2241\,
            I => \shift_regZ0Z_89\
        );

    \I__366\ : InMux
    port map (
            O => \N__2238\,
            I => \N__2235\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2235\,
            I => \shift_regZ0Z_54\
        );

    \I__364\ : InMux
    port map (
            O => \N__2232\,
            I => \N__2229\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2229\,
            I => \shift_regZ0Z_55\
        );

    \I__362\ : InMux
    port map (
            O => \N__2226\,
            I => \N__2223\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2223\,
            I => \shift_regZ0Z_56\
        );

    \I__360\ : InMux
    port map (
            O => \N__2220\,
            I => \N__2217\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2217\,
            I => \shift_regZ0Z_57\
        );

    \I__358\ : InMux
    port map (
            O => \N__2214\,
            I => \N__2211\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2211\,
            I => \shift_regZ0Z_58\
        );

    \I__356\ : InMux
    port map (
            O => \N__2208\,
            I => \N__2205\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2205\,
            I => \shift_regZ0Z_59\
        );

    \I__354\ : InMux
    port map (
            O => \N__2202\,
            I => \N__2199\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2199\,
            I => \N__2196\
        );

    \I__352\ : Odrv12
    port map (
            O => \N__2196\,
            I => \SPI_SDI_c\
        );

    \I__351\ : InMux
    port map (
            O => \N__2193\,
            I => \N__2190\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2190\,
            I => \shift_regZ0Z_0\
        );

    \I__349\ : InMux
    port map (
            O => \N__2187\,
            I => \N__2184\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2184\,
            I => \shift_regZ0Z_1\
        );

    \I__347\ : InMux
    port map (
            O => \N__2181\,
            I => \N__2178\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2178\,
            I => \shift_regZ0Z_2\
        );

    \I__345\ : InMux
    port map (
            O => \N__2175\,
            I => \N__2172\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__2172\,
            I => \shift_regZ0Z_61\
        );

    \I__343\ : InMux
    port map (
            O => \N__2169\,
            I => \N__2166\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2166\,
            I => \shift_regZ0Z_62\
        );

    \I__341\ : InMux
    port map (
            O => \N__2163\,
            I => \N__2160\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2160\,
            I => \shift_regZ0Z_63\
        );

    \I__339\ : InMux
    port map (
            O => \N__2157\,
            I => \N__2154\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2154\,
            I => \shift_regZ0Z_64\
        );

    \I__337\ : InMux
    port map (
            O => \N__2151\,
            I => \N__2148\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2148\,
            I => \shift_regZ0Z_65\
        );

    \I__335\ : InMux
    port map (
            O => \N__2145\,
            I => \N__2142\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2142\,
            I => \shift_regZ0Z_66\
        );

    \I__333\ : InMux
    port map (
            O => \N__2139\,
            I => \N__2136\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2136\,
            I => \shift_regZ0Z_51\
        );

    \I__331\ : InMux
    port map (
            O => \N__2133\,
            I => \N__2130\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2130\,
            I => \shift_regZ0Z_52\
        );

    \I__329\ : InMux
    port map (
            O => \N__2127\,
            I => \N__2124\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2124\,
            I => \shift_regZ0Z_53\
        );

    \I__327\ : InMux
    port map (
            O => \N__2121\,
            I => \N__2118\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2118\,
            I => \shift_regZ0Z_10\
        );

    \I__325\ : InMux
    port map (
            O => \N__2115\,
            I => \N__2112\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2112\,
            I => \shift_regZ0Z_11\
        );

    \I__323\ : InMux
    port map (
            O => \N__2109\,
            I => \N__2106\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2106\,
            I => \shift_regZ0Z_12\
        );

    \I__321\ : InMux
    port map (
            O => \N__2103\,
            I => \N__2100\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2100\,
            I => \shift_regZ0Z_13\
        );

    \I__319\ : InMux
    port map (
            O => \N__2097\,
            I => \N__2094\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2094\,
            I => \shift_regZ0Z_14\
        );

    \I__317\ : InMux
    port map (
            O => \N__2091\,
            I => \N__2088\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2088\,
            I => \shift_regZ0Z_15\
        );

    \I__315\ : InMux
    port map (
            O => \N__2085\,
            I => \N__2082\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2082\,
            I => \shift_regZ0Z_16\
        );

    \I__313\ : InMux
    port map (
            O => \N__2079\,
            I => \N__2076\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2076\,
            I => \shift_regZ0Z_17\
        );

    \I__311\ : InMux
    port map (
            O => \N__2073\,
            I => \N__2070\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2070\,
            I => \shift_regZ0Z_60\
        );

    \I__309\ : InMux
    port map (
            O => \N__2067\,
            I => \N__2064\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2064\,
            I => \shift_regZ0Z_6\
        );

    \I__307\ : InMux
    port map (
            O => \N__2061\,
            I => \N__2058\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2058\,
            I => \shift_regZ0Z_91\
        );

    \I__305\ : InMux
    port map (
            O => \N__2055\,
            I => \N__2052\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2052\,
            I => \shift_regZ0Z_92\
        );

    \I__303\ : InMux
    port map (
            O => \N__2049\,
            I => \N__2046\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2046\,
            I => \shift_regZ0Z_93\
        );

    \I__301\ : InMux
    port map (
            O => \N__2043\,
            I => \N__2040\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2040\,
            I => \shift_regZ0Z_94\
        );

    \I__299\ : InMux
    port map (
            O => \N__2037\,
            I => \N__2034\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2034\,
            I => \shift_regZ0Z_95\
        );

    \I__297\ : InMux
    port map (
            O => \N__2031\,
            I => \N__2028\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2028\,
            I => \shift_regZ0Z_7\
        );

    \I__295\ : InMux
    port map (
            O => \N__2025\,
            I => \N__2022\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2022\,
            I => \shift_regZ0Z_8\
        );

    \I__293\ : InMux
    port map (
            O => \N__2019\,
            I => \N__2016\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2016\,
            I => \shift_regZ0Z_9\
        );

    \I__291\ : InMux
    port map (
            O => \N__2013\,
            I => \N__2010\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2010\,
            I => \shift_regZ0Z_45\
        );

    \I__289\ : InMux
    port map (
            O => \N__2007\,
            I => \N__2004\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2004\,
            I => \shift_regZ0Z_46\
        );

    \I__287\ : InMux
    port map (
            O => \N__2001\,
            I => \N__1998\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__1998\,
            I => \shift_regZ0Z_47\
        );

    \I__285\ : InMux
    port map (
            O => \N__1995\,
            I => \N__1992\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__1992\,
            I => \shift_regZ0Z_48\
        );

    \I__283\ : InMux
    port map (
            O => \N__1989\,
            I => \N__1986\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__1986\,
            I => \shift_regZ0Z_49\
        );

    \I__281\ : InMux
    port map (
            O => \N__1983\,
            I => \N__1980\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__1980\,
            I => \shift_regZ0Z_50\
        );

    \I__279\ : InMux
    port map (
            O => \N__1977\,
            I => \N__1974\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__1974\,
            I => \shift_regZ0Z_96\
        );

    \I__277\ : InMux
    port map (
            O => \N__1971\,
            I => \N__1968\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__1968\,
            I => \shift_regZ0Z_97\
        );

    \I__275\ : InMux
    port map (
            O => \N__1965\,
            I => \N__1962\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__1962\,
            I => \shift_regZ0Z_108\
        );

    \I__273\ : CascadeMux
    port map (
            O => \N__1959\,
            I => \N__1956\
        );

    \I__272\ : InMux
    port map (
            O => \N__1956\,
            I => \N__1953\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__1953\,
            I => \shift_regZ0Z_109\
        );

    \I__270\ : InMux
    port map (
            O => \N__1950\,
            I => \N__1947\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__1947\,
            I => \shift_regZ0Z_103\
        );

    \I__268\ : InMux
    port map (
            O => \N__1944\,
            I => \N__1941\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__1941\,
            I => \shift_regZ0Z_104\
        );

    \I__266\ : InMux
    port map (
            O => \N__1938\,
            I => \N__1935\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__1935\,
            I => \shift_regZ0Z_105\
        );

    \I__264\ : InMux
    port map (
            O => \N__1932\,
            I => \N__1929\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__1929\,
            I => \shift_regZ0Z_106\
        );

    \I__262\ : InMux
    port map (
            O => \N__1926\,
            I => \N__1923\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__1923\,
            I => \shift_regZ0Z_107\
        );

    \I__260\ : InMux
    port map (
            O => \N__1920\,
            I => \N__1917\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__1917\,
            I => \shift_regZ0Z_18\
        );

    \I__258\ : InMux
    port map (
            O => \N__1914\,
            I => \N__1911\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__1911\,
            I => \shift_regZ0Z_19\
        );

    \I__256\ : InMux
    port map (
            O => \N__1908\,
            I => \N__1905\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__1905\,
            I => \shift_regZ0Z_43\
        );

    \I__254\ : InMux
    port map (
            O => \N__1902\,
            I => \N__1899\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__1899\,
            I => \shift_regZ0Z_44\
        );

    \I__252\ : InMux
    port map (
            O => \N__1896\,
            I => \N__1893\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__1893\,
            I => \shift_regZ0Z_100\
        );

    \I__250\ : InMux
    port map (
            O => \N__1890\,
            I => \N__1887\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1887\,
            I => \shift_regZ0Z_114\
        );

    \I__248\ : InMux
    port map (
            O => \N__1884\,
            I => \N__1881\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__1881\,
            I => \shift_regZ0Z_101\
        );

    \I__246\ : InMux
    port map (
            O => \N__1878\,
            I => \N__1875\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__1875\,
            I => \shift_regZ0Z_102\
        );

    \I__244\ : InMux
    port map (
            O => \N__1872\,
            I => \N__1869\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__1869\,
            I => \shift_regZ0Z_110\
        );

    \I__242\ : InMux
    port map (
            O => \N__1866\,
            I => \N__1863\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__1863\,
            I => \shift_regZ0Z_111\
        );

    \I__240\ : InMux
    port map (
            O => \N__1860\,
            I => \N__1857\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__1857\,
            I => \shift_regZ0Z_112\
        );

    \I__238\ : InMux
    port map (
            O => \N__1854\,
            I => \N__1851\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__1851\,
            I => \shift_regZ0Z_113\
        );

    \I__236\ : InMux
    port map (
            O => \N__1848\,
            I => \N__1845\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1845\,
            I => \shift_regZ0Z_37\
        );

    \I__234\ : InMux
    port map (
            O => \N__1842\,
            I => \N__1839\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__1839\,
            I => \shift_regZ0Z_38\
        );

    \I__232\ : InMux
    port map (
            O => \N__1836\,
            I => \N__1833\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__1833\,
            I => \shift_regZ0Z_39\
        );

    \I__230\ : InMux
    port map (
            O => \N__1830\,
            I => \N__1827\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__1827\,
            I => \shift_regZ0Z_40\
        );

    \I__228\ : InMux
    port map (
            O => \N__1824\,
            I => \N__1821\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__1821\,
            I => \shift_regZ0Z_41\
        );

    \I__226\ : InMux
    port map (
            O => \N__1818\,
            I => \N__1815\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__1815\,
            I => \shift_regZ0Z_42\
        );

    \I__224\ : InMux
    port map (
            O => \N__1812\,
            I => \N__1809\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__1809\,
            I => \shift_regZ0Z_98\
        );

    \I__222\ : InMux
    port map (
            O => \N__1806\,
            I => \N__1803\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1803\,
            I => \shift_regZ0Z_99\
        );

    \I__220\ : InMux
    port map (
            O => \N__1800\,
            I => \N__1797\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__1797\,
            I => \shift_regZ0Z_28\
        );

    \I__218\ : InMux
    port map (
            O => \N__1794\,
            I => \N__1791\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__1791\,
            I => \shift_regZ0Z_29\
        );

    \I__216\ : InMux
    port map (
            O => \N__1788\,
            I => \N__1785\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__1785\,
            I => \shift_regZ0Z_30\
        );

    \I__214\ : InMux
    port map (
            O => \N__1782\,
            I => \N__1779\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__1779\,
            I => \shift_regZ0Z_31\
        );

    \I__212\ : InMux
    port map (
            O => \N__1776\,
            I => \N__1773\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__1773\,
            I => \shift_regZ0Z_32\
        );

    \I__210\ : InMux
    port map (
            O => \N__1770\,
            I => \N__1767\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__1767\,
            I => \shift_regZ0Z_33\
        );

    \I__208\ : InMux
    port map (
            O => \N__1764\,
            I => \N__1761\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__1761\,
            I => \shift_regZ0Z_34\
        );

    \I__206\ : InMux
    port map (
            O => \N__1758\,
            I => \N__1755\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__1755\,
            I => \shift_regZ0Z_35\
        );

    \I__204\ : InMux
    port map (
            O => \N__1752\,
            I => \N__1749\
        );

    \I__203\ : LocalMux
    port map (
            O => \N__1749\,
            I => \shift_regZ0Z_36\
        );

    \I__202\ : InMux
    port map (
            O => \N__1746\,
            I => \N__1743\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__1743\,
            I => \shift_regZ0Z_115\
        );

    \I__200\ : InMux
    port map (
            O => \N__1740\,
            I => \N__1737\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__1737\,
            I => \shift_regZ0Z_20\
        );

    \I__198\ : InMux
    port map (
            O => \N__1734\,
            I => \N__1731\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__1731\,
            I => \shift_regZ0Z_21\
        );

    \I__196\ : InMux
    port map (
            O => \N__1728\,
            I => \N__1725\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1725\,
            I => \shift_regZ0Z_22\
        );

    \I__194\ : InMux
    port map (
            O => \N__1722\,
            I => \N__1719\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__1719\,
            I => \shift_regZ0Z_23\
        );

    \I__192\ : InMux
    port map (
            O => \N__1716\,
            I => \N__1713\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__1713\,
            I => \shift_regZ0Z_24\
        );

    \I__190\ : InMux
    port map (
            O => \N__1710\,
            I => \N__1707\
        );

    \I__189\ : LocalMux
    port map (
            O => \N__1707\,
            I => \shift_regZ0Z_25\
        );

    \I__188\ : InMux
    port map (
            O => \N__1704\,
            I => \N__1701\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__1701\,
            I => \shift_regZ0Z_26\
        );

    \I__186\ : InMux
    port map (
            O => \N__1698\,
            I => \N__1695\
        );

    \I__185\ : LocalMux
    port map (
            O => \N__1695\,
            I => \shift_regZ0Z_27\
        );

    \I__184\ : IoInMux
    port map (
            O => \N__1692\,
            I => \N__1689\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__1689\,
            I => \N__1686\
        );

    \I__182\ : Span4Mux_s2_v
    port map (
            O => \N__1686\,
            I => \N__1683\
        );

    \I__181\ : Odrv4
    port map (
            O => \N__1683\,
            I => \SPI_SDO_c\
        );

    \I__180\ : InMux
    port map (
            O => \N__1680\,
            I => \N__1677\
        );

    \I__179\ : LocalMux
    port map (
            O => \N__1677\,
            I => \shift_regZ0Z_119\
        );

    \I__178\ : InMux
    port map (
            O => \N__1674\,
            I => \N__1671\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1671\,
            I => \shift_regZ0Z_118\
        );

    \I__176\ : InMux
    port map (
            O => \N__1668\,
            I => \N__1665\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__1665\,
            I => \shift_regZ0Z_117\
        );

    \I__174\ : InMux
    port map (
            O => \N__1662\,
            I => \N__1659\
        );

    \I__173\ : LocalMux
    port map (
            O => \N__1659\,
            I => \shift_regZ0Z_116\
        );

    \I__172\ : ClkMux
    port map (
            O => \N__1656\,
            I => \N__1605\
        );

    \I__171\ : ClkMux
    port map (
            O => \N__1655\,
            I => \N__1605\
        );

    \I__170\ : ClkMux
    port map (
            O => \N__1654\,
            I => \N__1605\
        );

    \I__169\ : ClkMux
    port map (
            O => \N__1653\,
            I => \N__1605\
        );

    \I__168\ : ClkMux
    port map (
            O => \N__1652\,
            I => \N__1605\
        );

    \I__167\ : ClkMux
    port map (
            O => \N__1651\,
            I => \N__1605\
        );

    \I__166\ : ClkMux
    port map (
            O => \N__1650\,
            I => \N__1605\
        );

    \I__165\ : ClkMux
    port map (
            O => \N__1649\,
            I => \N__1605\
        );

    \I__164\ : ClkMux
    port map (
            O => \N__1648\,
            I => \N__1605\
        );

    \I__163\ : ClkMux
    port map (
            O => \N__1647\,
            I => \N__1605\
        );

    \I__162\ : ClkMux
    port map (
            O => \N__1646\,
            I => \N__1605\
        );

    \I__161\ : ClkMux
    port map (
            O => \N__1645\,
            I => \N__1605\
        );

    \I__160\ : ClkMux
    port map (
            O => \N__1644\,
            I => \N__1605\
        );

    \I__159\ : ClkMux
    port map (
            O => \N__1643\,
            I => \N__1605\
        );

    \I__158\ : ClkMux
    port map (
            O => \N__1642\,
            I => \N__1605\
        );

    \I__157\ : ClkMux
    port map (
            O => \N__1641\,
            I => \N__1605\
        );

    \I__156\ : ClkMux
    port map (
            O => \N__1640\,
            I => \N__1605\
        );

    \I__155\ : GlobalMux
    port map (
            O => \N__1605\,
            I => \N__1602\
        );

    \I__154\ : gio2CtrlBuf
    port map (
            O => \N__1602\,
            I => \SPI_SCK_c_g\
        );

    \I__153\ : IoInMux
    port map (
            O => \N__1599\,
            I => \N__1596\
        );

    \I__152\ : LocalMux
    port map (
            O => \N__1596\,
            I => \N__1593\
        );

    \I__151\ : Span4Mux_s1_h
    port map (
            O => \N__1593\,
            I => \N__1590\
        );

    \I__150\ : Span4Mux_h
    port map (
            O => \N__1590\,
            I => \N__1587\
        );

    \I__149\ : Odrv4
    port map (
            O => \N__1587\,
            I => \SPI_SCK_ibuf_gb_io_gb_input\
        );

    \INVshift_reg_68C\ : INV
    port map (
            O => \INVshift_reg_68C_net\,
            I => \N__1655\
        );

    \INVshift_reg_76C\ : INV
    port map (
            O => \INVshift_reg_76C_net\,
            I => \N__1647\
        );

    \INVshift_reg_90C\ : INV
    port map (
            O => \INVshift_reg_90C_net\,
            I => \N__1654\
        );

    \INVshift_reg_0C\ : INV
    port map (
            O => \INVshift_reg_0C_net\,
            I => \N__1656\
        );

    \INVshift_reg_52C\ : INV
    port map (
            O => \INVshift_reg_52C_net\,
            I => \N__1653\
        );

    \INVshift_reg_60C\ : INV
    port map (
            O => \INVshift_reg_60C_net\,
            I => \N__1651\
        );

    \INVshift_reg_10C\ : INV
    port map (
            O => \INVshift_reg_10C_net\,
            I => \N__1644\
        );

    \INVshift_reg_9C\ : INV
    port map (
            O => \INVshift_reg_9C_net\,
            I => \N__1650\
        );

    \INVshift_reg_96C\ : INV
    port map (
            O => \INVshift_reg_96C_net\,
            I => \N__1652\
        );

    \INVshift_reg_44C\ : INV
    port map (
            O => \INVshift_reg_44C_net\,
            I => \N__1649\
        );

    \INVshift_reg_108C\ : INV
    port map (
            O => \INVshift_reg_108C_net\,
            I => \N__1641\
        );

    \INVshift_reg_114C\ : INV
    port map (
            O => \INVshift_reg_114C_net\,
            I => \N__1646\
        );

    \INVshift_reg_98C\ : INV
    port map (
            O => \INVshift_reg_98C_net\,
            I => \N__1648\
        );

    \INVshift_reg_36C\ : INV
    port map (
            O => \INVshift_reg_36C_net\,
            I => \N__1645\
        );

    \INVshift_reg_28C\ : INV
    port map (
            O => \INVshift_reg_28C_net\,
            I => \N__1643\
        );

    \INVshift_reg_20C\ : INV
    port map (
            O => \INVshift_reg_20C_net\,
            I => \N__1640\
        );

    \INVSPI_SDOZ0C\ : INV
    port map (
            O => \INVSPI_SDOZ0C_net\,
            I => \N__1642\
        );

    \SPI_SCK_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1599\,
            GLOBALBUFFEROUTPUT => \SPI_SCK_c_g\
        );

    \SPI_SS_ibuf_RNIMF4D_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2370\,
            GLOBALBUFFEROUTPUT => \LED_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \SPI_SDOZ0_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1680\,
            lcout => \SPI_SDO_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVSPI_SDOZ0C_net\,
            ce => \N__2433\,
            sr => \_gnd_net_\
        );

    \shift_reg_119_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1674\,
            lcout => \shift_regZ0Z_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVSPI_SDOZ0C_net\,
            ce => \N__2433\,
            sr => \_gnd_net_\
        );

    \shift_reg_118_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1668\,
            lcout => \shift_regZ0Z_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVSPI_SDOZ0C_net\,
            ce => \N__2433\,
            sr => \_gnd_net_\
        );

    \shift_reg_117_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1662\,
            lcout => \shift_regZ0Z_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVSPI_SDOZ0C_net\,
            ce => \N__2433\,
            sr => \_gnd_net_\
        );

    \shift_reg_116_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1746\,
            lcout => \shift_regZ0Z_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVSPI_SDOZ0C_net\,
            ce => \N__2433\,
            sr => \_gnd_net_\
        );

    \shift_reg_115_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1890\,
            lcout => \shift_regZ0Z_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVSPI_SDOZ0C_net\,
            ce => \N__2433\,
            sr => \_gnd_net_\
        );

    \shift_reg_20_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1914\,
            lcout => \shift_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_20C_net\,
            ce => \N__2430\,
            sr => \_gnd_net_\
        );

    \shift_reg_21_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1740\,
            lcout => \shift_regZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_20C_net\,
            ce => \N__2430\,
            sr => \_gnd_net_\
        );

    \shift_reg_22_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1734\,
            lcout => \shift_regZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_20C_net\,
            ce => \N__2430\,
            sr => \_gnd_net_\
        );

    \shift_reg_23_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1728\,
            lcout => \shift_regZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_20C_net\,
            ce => \N__2430\,
            sr => \_gnd_net_\
        );

    \shift_reg_24_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1722\,
            lcout => \shift_regZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_20C_net\,
            ce => \N__2430\,
            sr => \_gnd_net_\
        );

    \shift_reg_25_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1716\,
            lcout => \shift_regZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_20C_net\,
            ce => \N__2430\,
            sr => \_gnd_net_\
        );

    \shift_reg_26_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1710\,
            lcout => \shift_regZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_20C_net\,
            ce => \N__2430\,
            sr => \_gnd_net_\
        );

    \shift_reg_27_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1704\,
            lcout => \shift_regZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_20C_net\,
            ce => \N__2430\,
            sr => \_gnd_net_\
        );

    \shift_reg_28_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1698\,
            lcout => \shift_regZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_28C_net\,
            ce => \N__2429\,
            sr => \_gnd_net_\
        );

    \shift_reg_29_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1800\,
            lcout => \shift_regZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_28C_net\,
            ce => \N__2429\,
            sr => \_gnd_net_\
        );

    \shift_reg_30_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1794\,
            lcout => \shift_regZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_28C_net\,
            ce => \N__2429\,
            sr => \_gnd_net_\
        );

    \shift_reg_31_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1788\,
            lcout => \shift_regZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_28C_net\,
            ce => \N__2429\,
            sr => \_gnd_net_\
        );

    \shift_reg_32_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1782\,
            lcout => \shift_regZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_28C_net\,
            ce => \N__2429\,
            sr => \_gnd_net_\
        );

    \shift_reg_33_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1776\,
            lcout => \shift_regZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_28C_net\,
            ce => \N__2429\,
            sr => \_gnd_net_\
        );

    \shift_reg_34_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1770\,
            lcout => \shift_regZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_28C_net\,
            ce => \N__2429\,
            sr => \_gnd_net_\
        );

    \shift_reg_35_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1764\,
            lcout => \shift_regZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_28C_net\,
            ce => \N__2429\,
            sr => \_gnd_net_\
        );

    \shift_reg_36_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1758\,
            lcout => \shift_regZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_36C_net\,
            ce => \N__2431\,
            sr => \_gnd_net_\
        );

    \shift_reg_37_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1752\,
            lcout => \shift_regZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_36C_net\,
            ce => \N__2431\,
            sr => \_gnd_net_\
        );

    \shift_reg_38_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1848\,
            lcout => \shift_regZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_36C_net\,
            ce => \N__2431\,
            sr => \_gnd_net_\
        );

    \shift_reg_39_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1842\,
            lcout => \shift_regZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_36C_net\,
            ce => \N__2431\,
            sr => \_gnd_net_\
        );

    \shift_reg_40_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1836\,
            lcout => \shift_regZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_36C_net\,
            ce => \N__2431\,
            sr => \_gnd_net_\
        );

    \shift_reg_41_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1830\,
            lcout => \shift_regZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_36C_net\,
            ce => \N__2431\,
            sr => \_gnd_net_\
        );

    \shift_reg_42_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1824\,
            lcout => \shift_regZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_36C_net\,
            ce => \N__2431\,
            sr => \_gnd_net_\
        );

    \shift_reg_43_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1818\,
            lcout => \shift_regZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_36C_net\,
            ce => \N__2431\,
            sr => \_gnd_net_\
        );

    \shift_reg_98_LC_3_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__1971\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \shift_regZ0Z_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_98C_net\,
            ce => \N__2440\,
            sr => \_gnd_net_\
        );

    \shift_reg_99_LC_3_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1812\,
            lcout => \shift_regZ0Z_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_98C_net\,
            ce => \N__2440\,
            sr => \_gnd_net_\
        );

    \shift_reg_100_LC_3_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1806\,
            lcout => \shift_regZ0Z_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_98C_net\,
            ce => \N__2440\,
            sr => \_gnd_net_\
        );

    \shift_reg_101_LC_3_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1896\,
            lcout => \shift_regZ0Z_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_98C_net\,
            ce => \N__2440\,
            sr => \_gnd_net_\
        );

    \shift_reg_114_LC_3_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1854\,
            lcout => \shift_regZ0Z_114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_114C_net\,
            ce => \N__2437\,
            sr => \_gnd_net_\
        );

    \shift_reg_102_LC_3_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1884\,
            lcout => \shift_regZ0Z_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_114C_net\,
            ce => \N__2437\,
            sr => \_gnd_net_\
        );

    \shift_reg_103_LC_3_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1878\,
            lcout => \shift_regZ0Z_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_114C_net\,
            ce => \N__2437\,
            sr => \_gnd_net_\
        );

    \shift_reg_110_LC_3_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1959\,
            in3 => \_gnd_net_\,
            lcout => \shift_regZ0Z_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_114C_net\,
            ce => \N__2437\,
            sr => \_gnd_net_\
        );

    \shift_reg_111_LC_3_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1872\,
            lcout => \shift_regZ0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_114C_net\,
            ce => \N__2437\,
            sr => \_gnd_net_\
        );

    \shift_reg_112_LC_3_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1866\,
            lcout => \shift_regZ0Z_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_114C_net\,
            ce => \N__2437\,
            sr => \_gnd_net_\
        );

    \shift_reg_113_LC_3_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1860\,
            lcout => \shift_regZ0Z_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_114C_net\,
            ce => \N__2437\,
            sr => \_gnd_net_\
        );

    \shift_reg_108_LC_3_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1926\,
            lcout => \shift_regZ0Z_108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_108C_net\,
            ce => \N__2434\,
            sr => \_gnd_net_\
        );

    \shift_reg_109_LC_3_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1965\,
            lcout => \shift_regZ0Z_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_108C_net\,
            ce => \N__2434\,
            sr => \_gnd_net_\
        );

    \shift_reg_104_LC_3_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1950\,
            lcout => \shift_regZ0Z_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_108C_net\,
            ce => \N__2434\,
            sr => \_gnd_net_\
        );

    \shift_reg_105_LC_3_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1944\,
            lcout => \shift_regZ0Z_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_108C_net\,
            ce => \N__2434\,
            sr => \_gnd_net_\
        );

    \shift_reg_106_LC_3_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1938\,
            lcout => \shift_regZ0Z_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_108C_net\,
            ce => \N__2434\,
            sr => \_gnd_net_\
        );

    \shift_reg_107_LC_3_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1932\,
            lcout => \shift_regZ0Z_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_108C_net\,
            ce => \N__2434\,
            sr => \_gnd_net_\
        );

    \shift_reg_18_LC_3_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2079\,
            lcout => \shift_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_108C_net\,
            ce => \N__2434\,
            sr => \_gnd_net_\
        );

    \shift_reg_19_LC_3_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1920\,
            lcout => \shift_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_108C_net\,
            ce => \N__2434\,
            sr => \_gnd_net_\
        );

    \shift_reg_44_LC_3_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1908\,
            lcout => \shift_regZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_44C_net\,
            ce => \N__2435\,
            sr => \_gnd_net_\
        );

    \shift_reg_45_LC_3_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1902\,
            lcout => \shift_regZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_44C_net\,
            ce => \N__2435\,
            sr => \_gnd_net_\
        );

    \shift_reg_46_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2013\,
            lcout => \shift_regZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_44C_net\,
            ce => \N__2435\,
            sr => \_gnd_net_\
        );

    \shift_reg_47_LC_3_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2007\,
            lcout => \shift_regZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_44C_net\,
            ce => \N__2435\,
            sr => \_gnd_net_\
        );

    \shift_reg_48_LC_3_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2001\,
            lcout => \shift_regZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_44C_net\,
            ce => \N__2435\,
            sr => \_gnd_net_\
        );

    \shift_reg_49_LC_3_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1995\,
            lcout => \shift_regZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_44C_net\,
            ce => \N__2435\,
            sr => \_gnd_net_\
        );

    \shift_reg_50_LC_3_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1989\,
            lcout => \shift_regZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_44C_net\,
            ce => \N__2435\,
            sr => \_gnd_net_\
        );

    \shift_reg_51_LC_3_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1983\,
            lcout => \shift_regZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_44C_net\,
            ce => \N__2435\,
            sr => \_gnd_net_\
        );

    \shift_reg_96_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2037\,
            lcout => \shift_regZ0Z_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_96C_net\,
            ce => \N__2443\,
            sr => \_gnd_net_\
        );

    \shift_reg_97_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1977\,
            lcout => \shift_regZ0Z_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_96C_net\,
            ce => \N__2443\,
            sr => \_gnd_net_\
        );

    \shift_reg_6_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2286\,
            lcout => \shift_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_96C_net\,
            ce => \N__2443\,
            sr => \_gnd_net_\
        );

    \shift_reg_7_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2067\,
            lcout => \shift_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_96C_net\,
            ce => \N__2443\,
            sr => \_gnd_net_\
        );

    \shift_reg_9_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2025\,
            lcout => \shift_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_9C_net\,
            ce => \N__2441\,
            sr => \_gnd_net_\
        );

    \shift_reg_91_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2280\,
            lcout => \shift_regZ0Z_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_9C_net\,
            ce => \N__2441\,
            sr => \_gnd_net_\
        );

    \shift_reg_92_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2061\,
            lcout => \shift_regZ0Z_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_9C_net\,
            ce => \N__2441\,
            sr => \_gnd_net_\
        );

    \shift_reg_93_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2055\,
            lcout => \shift_regZ0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_9C_net\,
            ce => \N__2441\,
            sr => \_gnd_net_\
        );

    \shift_reg_94_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2049\,
            lcout => \shift_regZ0Z_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_9C_net\,
            ce => \N__2441\,
            sr => \_gnd_net_\
        );

    \shift_reg_95_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2043\,
            lcout => \shift_regZ0Z_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_9C_net\,
            ce => \N__2441\,
            sr => \_gnd_net_\
        );

    \shift_reg_8_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2031\,
            lcout => \shift_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_9C_net\,
            ce => \N__2441\,
            sr => \_gnd_net_\
        );

    \shift_reg_10_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2019\,
            lcout => \shift_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_10C_net\,
            ce => \N__2438\,
            sr => \_gnd_net_\
        );

    \shift_reg_11_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2121\,
            lcout => \shift_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_10C_net\,
            ce => \N__2438\,
            sr => \_gnd_net_\
        );

    \shift_reg_12_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2115\,
            lcout => \shift_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_10C_net\,
            ce => \N__2438\,
            sr => \_gnd_net_\
        );

    \shift_reg_13_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2109\,
            lcout => \shift_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_10C_net\,
            ce => \N__2438\,
            sr => \_gnd_net_\
        );

    \shift_reg_14_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2103\,
            lcout => \shift_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_10C_net\,
            ce => \N__2438\,
            sr => \_gnd_net_\
        );

    \shift_reg_15_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2097\,
            lcout => \shift_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_10C_net\,
            ce => \N__2438\,
            sr => \_gnd_net_\
        );

    \shift_reg_16_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2091\,
            lcout => \shift_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_10C_net\,
            ce => \N__2438\,
            sr => \_gnd_net_\
        );

    \shift_reg_17_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2085\,
            lcout => \shift_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_10C_net\,
            ce => \N__2438\,
            sr => \_gnd_net_\
        );

    \shift_reg_60_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2208\,
            lcout => \shift_regZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_60C_net\,
            ce => \N__2432\,
            sr => \_gnd_net_\
        );

    \shift_reg_61_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2073\,
            lcout => \shift_regZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_60C_net\,
            ce => \N__2432\,
            sr => \_gnd_net_\
        );

    \shift_reg_62_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2175\,
            lcout => \shift_regZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_60C_net\,
            ce => \N__2432\,
            sr => \_gnd_net_\
        );

    \shift_reg_63_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2169\,
            lcout => \shift_regZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_60C_net\,
            ce => \N__2432\,
            sr => \_gnd_net_\
        );

    \shift_reg_64_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2163\,
            lcout => \shift_regZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_60C_net\,
            ce => \N__2432\,
            sr => \_gnd_net_\
        );

    \shift_reg_65_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2157\,
            lcout => \shift_regZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_60C_net\,
            ce => \N__2432\,
            sr => \_gnd_net_\
        );

    \shift_reg_66_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2151\,
            lcout => \shift_regZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_60C_net\,
            ce => \N__2432\,
            sr => \_gnd_net_\
        );

    \shift_reg_67_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2145\,
            lcout => \shift_regZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_60C_net\,
            ce => \N__2432\,
            sr => \_gnd_net_\
        );

    \shift_reg_52_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2139\,
            lcout => \shift_regZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_52C_net\,
            ce => \N__2439\,
            sr => \_gnd_net_\
        );

    \shift_reg_53_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2133\,
            lcout => \shift_regZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_52C_net\,
            ce => \N__2439\,
            sr => \_gnd_net_\
        );

    \shift_reg_54_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2127\,
            lcout => \shift_regZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_52C_net\,
            ce => \N__2439\,
            sr => \_gnd_net_\
        );

    \shift_reg_55_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2238\,
            lcout => \shift_regZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_52C_net\,
            ce => \N__2439\,
            sr => \_gnd_net_\
        );

    \shift_reg_56_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2232\,
            lcout => \shift_regZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_52C_net\,
            ce => \N__2439\,
            sr => \_gnd_net_\
        );

    \shift_reg_57_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2226\,
            lcout => \shift_regZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_52C_net\,
            ce => \N__2439\,
            sr => \_gnd_net_\
        );

    \shift_reg_58_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2220\,
            lcout => \shift_regZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_52C_net\,
            ce => \N__2439\,
            sr => \_gnd_net_\
        );

    \shift_reg_59_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2214\,
            lcout => \shift_regZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_52C_net\,
            ce => \N__2439\,
            sr => \_gnd_net_\
        );

    \shift_reg_0_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2202\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \shift_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_0C_net\,
            ce => \N__2445\,
            sr => \_gnd_net_\
        );

    \shift_reg_1_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2193\,
            lcout => \shift_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_0C_net\,
            ce => \N__2445\,
            sr => \_gnd_net_\
        );

    \shift_reg_2_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2187\,
            lcout => \shift_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_0C_net\,
            ce => \N__2445\,
            sr => \_gnd_net_\
        );

    \shift_reg_3_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2181\,
            lcout => \shift_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_0C_net\,
            ce => \N__2445\,
            sr => \_gnd_net_\
        );

    \shift_reg_4_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2298\,
            lcout => \shift_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_0C_net\,
            ce => \N__2445\,
            sr => \_gnd_net_\
        );

    \shift_reg_5_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2292\,
            lcout => \shift_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_0C_net\,
            ce => \N__2445\,
            sr => \_gnd_net_\
        );

    \shift_reg_90_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2244\,
            lcout => \shift_regZ0Z_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_90C_net\,
            ce => \N__2444\,
            sr => \_gnd_net_\
        );

    \shift_reg_84_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2310\,
            lcout => \shift_regZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_90C_net\,
            ce => \N__2444\,
            sr => \_gnd_net_\
        );

    \shift_reg_85_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2274\,
            lcout => \shift_regZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_90C_net\,
            ce => \N__2444\,
            sr => \_gnd_net_\
        );

    \shift_reg_86_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2268\,
            lcout => \shift_regZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_90C_net\,
            ce => \N__2444\,
            sr => \_gnd_net_\
        );

    \shift_reg_87_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2262\,
            lcout => \shift_regZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_90C_net\,
            ce => \N__2444\,
            sr => \_gnd_net_\
        );

    \shift_reg_88_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2256\,
            lcout => \shift_regZ0Z_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_90C_net\,
            ce => \N__2444\,
            sr => \_gnd_net_\
        );

    \shift_reg_89_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2250\,
            lcout => \shift_regZ0Z_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_90C_net\,
            ce => \N__2444\,
            sr => \_gnd_net_\
        );

    \shift_reg_76_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2451\,
            lcout => \shift_regZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_76C_net\,
            ce => \N__2442\,
            sr => \_gnd_net_\
        );

    \shift_reg_77_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2352\,
            lcout => \shift_regZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_76C_net\,
            ce => \N__2442\,
            sr => \_gnd_net_\
        );

    \shift_reg_78_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2346\,
            lcout => \shift_regZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_76C_net\,
            ce => \N__2442\,
            sr => \_gnd_net_\
        );

    \shift_reg_79_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2340\,
            lcout => \shift_regZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_76C_net\,
            ce => \N__2442\,
            sr => \_gnd_net_\
        );

    \shift_reg_80_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2334\,
            lcout => \shift_regZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_76C_net\,
            ce => \N__2442\,
            sr => \_gnd_net_\
        );

    \shift_reg_81_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2328\,
            lcout => \shift_regZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_76C_net\,
            ce => \N__2442\,
            sr => \_gnd_net_\
        );

    \shift_reg_82_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2322\,
            lcout => \shift_regZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_76C_net\,
            ce => \N__2442\,
            sr => \_gnd_net_\
        );

    \shift_reg_83_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2316\,
            lcout => \shift_regZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_76C_net\,
            ce => \N__2442\,
            sr => \_gnd_net_\
        );

    \shift_reg_68_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2304\,
            lcout => \shift_regZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_68C_net\,
            ce => \N__2436\,
            sr => \_gnd_net_\
        );

    \shift_reg_69_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2493\,
            lcout => \shift_regZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_68C_net\,
            ce => \N__2436\,
            sr => \_gnd_net_\
        );

    \shift_reg_70_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2487\,
            lcout => \shift_regZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_68C_net\,
            ce => \N__2436\,
            sr => \_gnd_net_\
        );

    \shift_reg_71_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2481\,
            lcout => \shift_regZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_68C_net\,
            ce => \N__2436\,
            sr => \_gnd_net_\
        );

    \shift_reg_72_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2475\,
            lcout => \shift_regZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_68C_net\,
            ce => \N__2436\,
            sr => \_gnd_net_\
        );

    \shift_reg_73_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2469\,
            lcout => \shift_regZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_68C_net\,
            ce => \N__2436\,
            sr => \_gnd_net_\
        );

    \shift_reg_74_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2463\,
            lcout => \shift_regZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_68C_net\,
            ce => \N__2436\,
            sr => \_gnd_net_\
        );

    \shift_reg_75_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2457\,
            lcout => \shift_regZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVshift_reg_68C_net\,
            ce => \N__2436\,
            sr => \_gnd_net_\
        );

    \SPI_SS_ibuf_RNIMF4D_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2387\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LED_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
